module Decodificador_binario_gray_tb();
	logic A, B, C, D;
	logic [6:0] seven_segment_pins;
	
	Decodificador_binario_gray dut (
        .A(A), 
        .B(B), 
        .C(C), 
        .D(D), 
        .seven_segment_pins(seven_segment_pins)
    );

    
    initial begin
        $display("Tiempo | Binario | Gray | 7-seg");
        $display("--------------------------------");

        // Número 0 (0000)
        A=0; B=0; C=0; D=0;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);
					  

			// Número 1 (0001)
        A=0; B=0; C=0; D=1;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);
					  
			// Número 2 (0010)
        A=0; B=0; C=1; D=0;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);
					  
		  // Número 3 (0011)
        A=0; B=0; C=1; D=1;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);
					  
		  // Número 4 (0100)
        A=0; B=1; C=0; D=0;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 5 (0101)
        A=0; B=1; C=0; D=1;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);
					  
		  // Número 6 (0110)
        A=0; B=1; C=1; D=0; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 7 (0111)
        A=0; B=1; C=1; D=1; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 8 (1000)
        A=1; B=0; C=0; D=0; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 9 (1001)
        A=1; B=0; C=0; D=1; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 10 (1010)
        A=1; B=0; C=1; D=0; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 11 (1011)
        A=1; B=0; C=1; D=1; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 12 (1100)
        A=1; B=1; C=0; D=0; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 13 (1101)
        A=1; B=1; C=0; D=1; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);

        // Número 14 (1110)
        A=1; B=1; C=1; D=0; #10;
        $display("%4t | %b%b%b%b | %b | %b", $time, A, B, C, D, dut.dec_result, seven_segment_pins);


        // Número 15 (1111)
        A=1; B=1; C=1; D=1;
        #10;
        $display("%4t   | %b%b%b%b   | %b   | %b", 
                 $time, A, B, C, D, dut.dec_result, seven_segment_pins);

       
    end
endmodule
